module ysyx_23060236_idu(
	input  [31:0] in,
	output [9:0]  opcode_type,
	output [2:0]  funct3,
	output [6:0]  funct7,
	output [3:0]  rd,
	output [3:0]  rs1,
	output [3:0]  rs2,
	output [31:0] imm,
	output lsu_wen,
	output lsu_ren,
	output reg_wen,
	output csr_enable,
	output inst_fencei,
	output inst_ecall,
	output inst_mret,
	input  idu_valid);

	wire [5:0] Type;
	wire [6:0] opcode;
	assign opcode  = in[6:0];
	assign rs1     = in[18:15];
	assign rs2     = in[23:20];
	assign rd      = in[10:7];
	assign funct3  = in[14:12];
	assign funct7  = in[31:25];
	assign lsu_ren = (opcode_type[INST_LW]) & idu_valid;
	assign lsu_wen = (opcode_type[INST_SW]) & idu_valid;
	assign reg_wen = Type[TYPE_I] & ~((funct3 == 3'b0) & opcode_type[INST_CSR]) | Type[TYPE_U] | Type[TYPE_J] | Type[TYPE_R];
	assign csr_enable = (opcode_type[INST_CSR]) & (funct3 != 3'b0);

	assign inst_ecall  = (in == 32'h00000073);
	assign inst_mret   = (in == 32'h30200073);
	assign inst_fencei = (opcode == 7'b0001111);

	parameter TYPE_R = 0;
	parameter TYPE_I = 1;
	parameter TYPE_S = 2;
	parameter TYPE_B = 3;
	parameter TYPE_U = 4;
	parameter TYPE_J = 5; 

	parameter INST_LUI   = 0;
	parameter INST_AUIPC = 1;
	parameter INST_JAL   = 2;
	parameter INST_JALR  = 3;
	parameter INST_BEQ   = 4;
	parameter INST_LW    = 5;
	parameter INST_SW    = 6;
	parameter INST_ADDI  = 7;
	parameter INST_ADD   = 8;
	parameter INST_CSR   = 9;

	assign opcode_type[INST_LUI  ] = (opcode == 7'b0110111);
	assign opcode_type[INST_AUIPC] = (opcode == 7'b0010111);
	assign opcode_type[INST_JAL  ] = (opcode == 7'b1101111);
	assign opcode_type[INST_JALR ] = (opcode == 7'b1100111);
	assign opcode_type[INST_BEQ  ] = (opcode == 7'b1100011);
	assign opcode_type[INST_LW   ] = (opcode == 7'b0000011);
	assign opcode_type[INST_SW   ] = (opcode == 7'b0100011);
	assign opcode_type[INST_ADDI ] = (opcode == 7'b0010011);
	assign opcode_type[INST_ADD  ] = (opcode == 7'b0110011);
	assign opcode_type[INST_CSR  ] = (opcode == 7'b1110011);

	assign Type[TYPE_R] = opcode_type[INST_ADD];
	assign Type[TYPE_I] = opcode_type[INST_JALR] | opcode_type[INST_LW] | opcode_type[INST_ADDI] | opcode_type[INST_CSR];
	assign Type[TYPE_S] = opcode_type[INST_SW];
	assign Type[TYPE_B] = opcode_type[INST_BEQ];
	assign Type[TYPE_U] = opcode_type[INST_LUI] | opcode_type[INST_AUIPC];
	assign Type[TYPE_J] = opcode_type[INST_JAL];

	assign imm = (Type[TYPE_I]) ? {{20{in[31]}}, in[31:20]} :
	             (Type[TYPE_U]) ? {in[31:12], 12'b0} :
	             (Type[TYPE_S]) ? {{20{in[31]}}, in[31:25], in[11:7]} :
	             (Type[TYPE_J]) ? {{12{in[31]}}, in[19:12], in[20], in[30:21], 1'b0} :
	             (Type[TYPE_B]) ? {{20{in[31]}}, in[7], in[30:25], in[11:8], 1'b0} :
							 32'b0;

endmodule
