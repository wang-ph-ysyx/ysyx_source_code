module ysyx_23060236_ifu(
	input  clock,
	input  reset,

	output [31:0] ifu_araddr,
	output        ifu_arvalid,
	input         ifu_arready,
	input  [63:0] ifu_rdata,
	input  [1:0]  ifu_rresp,
	input         ifu_rvalid,
	output        ifu_rready,

	output [31:0] icache_araddr,
	output        icache_arvalid,
	input         icache_arready,
	input  [31:0] icache_rdata,
	input  [1:0]  icache_rresp,
	input         icache_rvalid,
	output        icache_rready,

	output        icache_awvalid,
	output [31:0] icache_awaddr,
	input         icache_awready,
	output [31:0] icache_wdata,
	output [7:0]  icache_wstrb,
	output        icache_wvalid,
	input         icache_wready,
	input  [1:0]  icache_bresp,
	input         icache_bvalid,
	output        icache_bready,


	input         wb_valid,
	input  [31:0] pc,
	output [31:0] inst,
	output        ifu_aligned,
	output        idu_valid
);

	wire [31:0] inst_tmp;
	wire [31:0] inst_icache_tmp;
	wire [31:0] inst_ifu_tmp;

	assign icache_rready = 1;
	assign icache_araddr = pc;
	assign icache_awaddr = pc;
	assign icache_wdata  = inst;
	assign icache_wstrb  = 8'hff;
	assign icache_bready = 1;
	assign ifu_rready    = 1;
	assign ifu_araddr    = pc;
	assign ifu_aligned   = (ifu_araddr >= 32'h0f000000) & (ifu_araddr < 32'h0f002000);
	assign inst_ifu_tmp  = ({32{~ifu_aligned}} & ifu_rdata[31:0] | {32{ifu_aligned}} & ({32{pc[2]}} & ifu_rdata[63:32] | {32{~pc[2]}} & ifu_rdata[31:0])) & {32{ifu_rvalid & ifu_rready}};
	assign inst_icache_tmp = icache_rdata & {32{icache_rvalid & icache_rready & ~icache_rresp[1]}};
	assign inst_tmp = inst_ifu_tmp | inst_icache_tmp;

	ysyx_23060236_Reg #(1, 0) reg_icache_arvalid(
		.clock(clock),
		.reset(reset),
		.din(icache_arvalid & ~icache_arready | ~icache_arvalid & wb_valid),
		.dout(icache_arvalid),
		.wen(1)
	);

	ysyx_23060236_Reg #(1, 0) reg_icache_awvalid(
		.clock(clock),
		.reset(reset),
		.din(icache_awvalid & ~icache_awready | ~icache_awvalid & icache_rvalid & icache_rready & icache_rresp[1]),
		.dout(icache_awvalid),
		.wen(1)
	);

	ysyx_23060236_Reg #(1, 0) reg_icache_wvalid(
		.clock(clock),
		.reset(reset),
		.din(icache_wvalid & ~icache_wready | ~icache_wvalid & ifu_rvalid & ifu_rready),
		.dout(icache_wvalid),
		.wen(1)
	);

	ysyx_23060236_Reg #(1, 1) reg_ifu_arvalid(
		.clock(clock),
		.reset(reset),
		.din(ifu_arvalid & ~ifu_arready | ~ifu_arvalid & (icache_rvalid & icache_rready & icache_rresp[1])),
		.dout(ifu_arvalid),
		.wen(1)
	);

	ysyx_23060236_Reg #(32, 0) reg_inst(
		.clock(clock),
		.reset(reset),
		.din(inst_tmp),
		.dout(inst),
		.wen(ifu_rvalid & ifu_rready | icache_rvalid & icache_rready & ~icache_rresp[1])
	);

	ysyx_23060236_Reg #(1, 0) reg_idu_valid(
		.clock(clock),
		.reset(reset),
		.din(~idu_valid & (icache_rvalid & icache_rready & ~icache_rresp[1] | icache_bvalid & icache_bready)),
		.dout(idu_valid),
		.wen(1)
	);

endmodule
