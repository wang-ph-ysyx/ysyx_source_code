`include "ysyx_23060236_defines.v"
module ysyx_23060236_lsu(
	input  clock,
	input  reset,

	output [31:0] lsu_araddr,
	output        lsu_arvalid,
	output [2:0]  lsu_arsize,
	input         lsu_arready,
	input  [31:0] lsu_rdata,
	input  [1:0]  lsu_rresp,
	input         lsu_rvalid,
	output        lsu_rready,

	output [31:0] lsu_awaddr,
	output        lsu_awvalid,
	output [2:0]  lsu_awsize,
	input         lsu_awready,
	output [31:0] lsu_wdata,
	output [3:0]  lsu_wstrb,
	output        lsu_wvalid,
	input         lsu_wready,
	input  [1:0]  lsu_bresp,
	input         lsu_bvalid,
	output        lsu_bready,

	input  [31:0] exu_val,
	input  [31:0] muldiv_val,
	input  [31:0] lsu_data,
	input  lsu_ren,
	input  lsu_wen,
	input  jump_wrong,
	input  [2:0]  funct3_reg,

	output reg [31:0] wb_val,

	input  inst_muldiv,
	input  muldiv_outvalid,
	input  exu_valid,
	input  exu_ready,
	output lsu_over,
	output wb_valid,

	input  time_intr,

	output [31:0] dcache_araddr,
	input  [31:0] dcache_rdata,
	input                 dcache_hit,  

	output [31:0] dcache_awaddr,
	output [31:0] dcache_wdata,
	output        dcache_wvalid,
	output        dirty_data,

	input             dcache_wdt,
	input  reg [25:0] dcache_reptag, //与dcache的tag位宽一致
	input  reg [31:0] dcache_repdata,

	output flush
);

	reg  [31:0] lsu_data_reg;
	wire [31:0] lsu_addr;
	wire [3:0]  wmask;
	wire handshake;

	assign handshake = exu_valid & exu_ready & ~time_intr;
	assign lsu_over = handshake & ~lsu_ren & ~lsu_wen & ~inst_muldiv | 
										lsu_rvalid & lsu_rready |	
										lsu_bvalid & lsu_bready | 
										muldiv_outvalid;
	assign lsu_addr = wb_val;
	assign wmask = (funct3_reg[1:0] == 2'b00) ? 4'h1 : 
								 (funct3_reg[1:0] == 2'b01) ? 4'h3 :
								 (funct3_reg[1:0] == 2'b10) ? 4'hf : 
								 4'b0;

	always @(posedge clock) begin
		if (handshake) begin
			wb_val          <= exu_val;
			lsu_data_reg    <= lsu_data;
		end
		else if (lsu_rvalid & lsu_rready) begin
			wb_val <= lsu_val_tmp;
		end
		else if (muldiv_outvalid) begin
			wb_val <= muldiv_val;
		end
	end

	ysyx_23060236_Reg #(1, 0) reg_wb_valid(
		.clock(clock),
		.reset(reset),
		.din(lsu_over),
		.dout(wb_valid),
		.wen(1)
	);

	wire [31:0] lsu_val_tmp;
	wire [31:0] lsu_val_shift;

	assign lsu_arsize = {1'b0, funct3_reg[1:0]};
	assign lsu_awsize = {1'b0, funct3_reg[1:0]};
	assign lsu_rready = 1;
	assign lsu_bready = 1;
	assign lsu_araddr = lsu_addr;
	assign lsu_awaddr = lsu_addr;
	assign lsu_wstrb  = wmask << lsu_awaddr[1:0];
	assign lsu_wdata  = lsu_data_reg << {lsu_awaddr[1:0], 3'b0};
	assign lsu_val_shift = lsu_rdata >> {lsu_araddr[1:0], 3'b0};

	assign lsu_val_tmp = (funct3_reg == 3'b000) ? (lsu_val_shift & 32'hff) | {{24{lsu_val_shift[7]}}, 8'h0} :     //lb  
                       (funct3_reg == 3'b001) ? (lsu_val_shift & 32'hffff) | {{16{lsu_val_shift[15]}}, 16'h0} : //lh
                       (funct3_reg == 3'b010) ? lsu_val_shift :                                                 //lw
                       (funct3_reg == 3'b100) ? lsu_val_shift & 32'hff :                                        //lbu
                       (funct3_reg == 3'b101) ? lsu_val_shift & 32'hffff :                                      //lhu
											 32'b0;

	ysyx_23060236_Reg #(1, 0) reg_lsu_arvalid(
		.clock(clock),
		.reset(reset),
		.din(lsu_arvalid & ~lsu_arready | ~lsu_arvalid & lsu_ren & handshake),
		.dout(lsu_arvalid),
		.wen(1)
	);

	ysyx_23060236_Reg #(1, 0) reg_lsu_awvalid(
		.clock(clock),
		.reset(reset),
		.din(lsu_awvalid & ~lsu_awready | ~lsu_awvalid & lsu_wen & handshake),
		.dout(lsu_awvalid),
		.wen(1)
	);

	ysyx_23060236_Reg #(1, 0) reg_lsu_wvalid(
		.clock(clock),
		.reset(reset),
		.din(lsu_wvalid & ~lsu_wready | ~lsu_wvalid & lsu_wen & handshake),
		.dout(lsu_wvalid),
		.wen(1)
	);

endmodule
