module ysyx_23060236_CSRFile #(DATA_WIDTH = 1) (
	input clock,
	input [11:0] imm,
	input [DATA_WIDTH-1:0] wdata,
	output [DATA_WIDTH-1:0] rdata,
	input enable,
	input inst_ecall,
	input [31:0] epc,
	input [31:0] cause,
	output [31:0] jump,
	input inst_mret,
	input valid
);

	wire [2:0] addr;
	reg [DATA_WIDTH-1:0] csr [5:0];//0:mepc  1:mcause  2:mstatus  3:mtvec  4:mvendorid  5:marchid

	ysyx_23060236_MuxKeyInternal #(6, 12, 3, 1) choose_addr(
		.out(addr),
		.key(imm),
		.default_out(3'b000),
		.lut({
			12'h341, 3'b000, //mepc
			12'h342, 3'b001, //mcause
			12'h300, 3'b010, //mstatus
			12'h305, 3'b011, //mtvec
			12'hf11, 3'b100, //mvendorid
			12'hf12, 3'b101  //marchid
		})
	);

	always @(posedge clock) begin
		if (valid) begin
			if (enable) begin
				csr[addr] <= wdata;
			end
			else if (inst_ecall) begin
				csr[0] <= epc + 4;
				csr[1] <= cause;
			end else begin
				csr[4] <= 32'h79737978;
				csr[5] <= 32'h015fdf0c;
			end
		end
	end

	assign rdata = {32{enable}} & csr[addr];
	assign jump = {32{inst_ecall}} & csr[3] | {32{inst_mret}} & csr[0];

endmodule
