module ysyx_23060236_lsu(
	input  clock,
	input  reset,

	output [31:0] lsu_araddr,
	output        lsu_arvalid,
	output [2:0]  lsu_arsize,
	input         lsu_arready,
	input  [63:0] lsu_rdata,
	input  [1:0]  lsu_rresp,
	input         lsu_rvalid,
	output        lsu_rready,

	output [31:0] lsu_awaddr,
	output        lsu_awvalid,
	output [2:0]  lsu_awsize,
	input         lsu_awready,
	output [63:0] lsu_wdata,
	output [7:0]  lsu_wstrb,
	output        lsu_wvalid,
	input         lsu_wready,
	input  [1:0]  lsu_bresp,
	input         lsu_bvalid,
	output        lsu_bready,

	input  [6:0]  opcode,
	input  [2:0]  funct3,
	input  [31:0] src1,
	input  [31:0] src2,
	input  [31:0] imm,
	input  [7:0]  wmask,
	input         wb_valid,
	input         lsu_ren,
	input         lsu_wen,
	output        lsu_aligned_64,
	output        lsu_aligned_32,
	output [31:0] lsu_val
);

	wire [31:0] lsu_val_raw;
	wire [31:0] lsu_val_tmp;
	wire [31:0] lsu_val_shift;
	wire [31:0] lsu_rdata_32;

	assign lsu_arsize = {1'b0, funct3[1:0]};
	assign lsu_awsize = {1'b0, funct3[1:0]};

	ysyx_23060236_MuxKeyInternal #(5, 3, 32, 1) caculate_lsu_val_tmp(
		.out(lsu_val_tmp),
		.key(funct3),
		.default_out(32'b0),
		.lut({
			3'b000, (lsu_val_raw & 32'hff) | {{24{lsu_val_raw[7]}}, 8'h0},      //lb
			3'b001, (lsu_val_raw & 32'hffff) | {{16{lsu_val_raw[15]}}, 16'h0},  //lh
			3'b010, lsu_val_raw,                                                //lw
			3'b100, lsu_val_raw & 32'hff,                                       //lbu
			3'b101, lsu_val_raw & 32'hffff                                      //lhu
		})
	);

	ysyx_23060236_MuxKeyInternal #(4, 2, 32, 1) calculate_lsu_val_shift(
		.out(lsu_val_shift),
		.key(lsu_araddr[1:0]),
		.default_out(32'b0),
		.lut({
			2'b00, lsu_rdata_32[31:0],
			2'b01, {8'b0,  lsu_rdata_32[31:8]},
			2'b10, {16'b0, lsu_rdata_32[31:16]},
			2'b11, {24'b0, lsu_rdata_32[31:24]}
		})
	);

	ysyx_23060236_MuxKeyInternal #(8, 3, 8, 1) calculate_lsu_wstrb(
		.out(lsu_wstrb),
		.key(lsu_awaddr[2:0]),
		.default_out(8'b0),
		.lut({
			3'b000, wmask,
			3'b001, {wmask[6:0], 1'b0},
			3'b010, {wmask[5:0], 2'b0},
			3'b011, {wmask[4:0], 3'b0},
			3'b100, {wmask[3:0], 4'b0},
			3'b101, {wmask[2:0], 5'b0},
			3'b110, {wmask[1:0], 6'b0},
			3'b111, {wmask[0:0], 7'b0}
		})
	);

	assign lsu_wdata = {32'b0, src2} << {lsu_awaddr[2:0], 3'b0};

	ysyx_23060236_Reg #(32, 0) reg_lsu_val(
		.clock(clock),
		.reset(reset),
		.din(lsu_val_tmp & {32{~wb_valid}}),
		.dout(lsu_val),
		.wen(lsu_rvalid & lsu_rready | wb_valid)
	);

	ysyx_23060236_Reg #(1, 0) reg_lsu_arvalid(
		.clock(clock),
		.reset(reset),
		.din(lsu_arvalid & ~lsu_arready | ~lsu_arvalid & lsu_ren),
		.dout(lsu_arvalid),
		.wen(1)
	);

	ysyx_23060236_Reg #(1, 0) reg_lsu_awvalid(
		.clock(clock),
		.reset(reset),
		.din(lsu_awvalid & ~lsu_awready | ~lsu_awvalid & lsu_wen),
		.dout(lsu_awvalid),
		.wen(1)
	);

	ysyx_23060236_Reg #(1, 0) reg_lsu_wvalid(
		.clock(clock),
		.reset(reset),
		.din(lsu_wvalid & ~lsu_wready | ~lsu_wvalid & lsu_wen),
		.dout(lsu_wvalid),
		.wen(1)
	);

	assign lsu_rready = 1;
	assign lsu_bready = 1;
	assign lsu_araddr = src1 + imm;
	assign lsu_awaddr = src1 + imm;
	assign lsu_aligned_64 = (lsu_araddr >= 32'h0f000000) & (lsu_araddr < 32'h0f002000);
	assign lsu_aligned_32 = (lsu_araddr >= 32'h80000000) & (lsu_araddr < 32'hc0000000);
	assign lsu_rdata_32 = (lsu_aligned_64 & lsu_araddr[2]) ? lsu_rdata[63:32] : lsu_rdata[31:0];
	assign lsu_val_raw = (lsu_aligned_64 | lsu_aligned_32) ? lsu_val_shift : lsu_rdata_32;

endmodule
