module ysyx_23060236_CSRFile #(DATA_WIDTH = 32) (
	input  clock,
	input  reset,
	input  [11:0] read_imm,
	input  [11:0] write_imm,
	input  [DATA_WIDTH-1:0] wdata,
	output [DATA_WIDTH-1:0] rdata,
	input  enable,
	input  inst_ecall,
	input  inst_ecall_write,
	input  inst_mret,
	input  [31:0] epc,
	output [31:0] jump,
	output        jump_en,
	input  valid
);

	reg [DATA_WIDTH-1:0] mepc   ;
	reg [DATA_WIDTH-1:0] mcause ;
	reg [DATA_WIDTH-1:0] mstatus;
	reg [DATA_WIDTH-1:0] mtvec  ;

	always @(posedge clock) begin
		if (reset) begin
			mstatus <= 32'h1800;
		end
		else if (valid) begin
			if (enable) begin
				if (write_imm == 12'h341) mepc    <= wdata;
				if (write_imm == 12'h342) mcause  <= wdata;
				if (write_imm == 12'h300) mstatus <= wdata;
				if (write_imm == 12'h305) mtvec   <= wdata;
			end
			else if (inst_ecall_write) begin
				mepc   <= epc;
				mcause <= 32'd11;
			end
		end
	end

	assign rdata = (read_imm == 12'h341) ? mepc    :
                 (read_imm == 12'h342) ? mcause  :
                 (read_imm == 12'h300) ? mstatus :
                 (read_imm == 12'h305) ? mtvec   :
                 (read_imm == 12'hf11) ? 32'h79737978 :
                 (read_imm == 12'hf12) ? 32'h015fdf0c :
								 32'b0;

	assign jump = {32{inst_ecall}} & mtvec | {32{inst_mret}} & mepc;
	assign jump_en = inst_ecall | inst_mret;

endmodule
