module idu(
	input [31:0] in,
	output [6:0] opcode,
	output [2:0] funct3,
	output [6:0] funct7,
	output [4:0] rd,
	output [4:0] rs1,
	output [4:0] rs2,
	output [31:0] imm,
	output [2:0] Type);

	assign opcode = in[6:0];
	assign rs1 = in[19:15];
	assign rs2 = in[24:20];
	assign rd = in[11:7];
	assign funct3 = in[14:12];

	parameter TYPE_R = 3'd0, TYPE_I = 3'd1, TYPE_S = 3'd2, TYPE_B = 3'd3, TYPE_U = 3'd4, TYPE_J = 3'd5; 

	MuxKeyInternal #(1, 7, 3, 0) choose_type(
		.out(Type),
		.key(opcode),
		.default_out(3'b0),
		.lut({
			7'b0010011, TYPE_I
		})
	);

	MuxKeyInternal #(1, 3, 32, 0) choose_imm(
		.out(imm),
		.key(Type),
		.default_out(32'b0),
		.lut({
			TYPE_I, {20'b0, in[31:20]}
		})
	);

endmodule
