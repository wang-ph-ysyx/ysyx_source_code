module npc(
	input  clock,
	input  reset,
);

  ysyx_23060236 cpu (	
    .clock                   (clock),
    .reset                   (reset),
    .io_interrupt            (1'h0),
    .io_master_awready      (auto_master_out_awready),
    .io_master_awvalid      (auto_master_out_awvalid),
    .io_master_awid    (auto_master_out_awid),
    .io_master_awaddr  (auto_master_out_awaddr),
    .io_master_awlen   (auto_master_out_awlen),
    .io_master_awsize  (auto_master_out_awsize),
    .io_master_awburst (auto_master_out_awburst),
    .io_master_wready       (auto_master_out_wready),
    .io_master_wvalid       (auto_master_out_wvalid),
    .io_master_wdata   (auto_master_out_wdata),
    .io_master_wstrb   (auto_master_out_wstrb),
    .io_master_wlast   (auto_master_out_wlast),
    .io_master_bready       (auto_master_out_bready),
    .io_master_bvalid       (auto_master_out_bvalid),
    .io_master_bid     (auto_master_out_bid),
    .io_master_bresp   (auto_master_out_bresp),
    .io_master_arready      (auto_master_out_arready),
    .io_master_arvalid      (auto_master_out_arvalid),
    .io_master_arid    (auto_master_out_arid),
    .io_master_araddr  (auto_master_out_araddr),
    .io_master_arlen   (auto_master_out_arlen),
    .io_master_arsize  (auto_master_out_arsize),
    .io_master_arburst (auto_master_out_arburst),
    .io_master_rready       (auto_master_out_rready),
    .io_master_rvalid       (auto_master_out_rvalid),
    .io_master_rid     (auto_master_out_rid),
    .io_master_rdata   (auto_master_out_rdata),
    .io_master_rresp   (auto_master_out_rresp),
    .io_master_rlast   (auto_master_out_rlast),
    .io_slave_awready       (/* unused */),
    .io_slave_awvalid       (1'h0),	
    .io_slave_awid     (4'h0),	
    .io_slave_awaddr   (32'h0),	
    .io_slave_awlen    (8'h0),	
    .io_slave_awsize   (3'h0),	
    .io_slave_awburst  (2'h0),	
    .io_slave_wready        (/* unused */),
    .io_slave_wvalid        (1'h0),	
    .io_slave_wdata    (32'h0),	
    .io_slave_wstrb    (4'h0),	
    .io_slave_wlast    (1'h0),	
    .io_slave_bready        (1'h0),	
    .io_slave_bvalid        (/* unused */),
    .io_slave_bid      (/* unused */),
    .io_slave_bresp    (/* unused */),
    .io_slave_arready       (/* unused */),
	);

endmodule
